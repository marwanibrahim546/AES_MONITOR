class AES_monitor_before extends uvm_monitor;

	`uvm_component_utils(AES_monitor_before)






endclass : AES_monitor_before

////////////////////////////////////////////////////////////////////

class AES_monitor_after extends uvm_monitor;

	`uvm_component_utils(AES_monitor_after)






endclass : AES_monitor_after